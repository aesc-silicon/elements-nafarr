module USRMCLK (
	input USRMCLKI,
	input USRMCLKTS
);

endmodule
