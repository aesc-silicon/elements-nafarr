// SPDX-FileCopyrightText: 2025 aesc silicon
//
// SPDX-License-Identifier: CERN-OHL-W-2.0

module USRMCLK (
	input USRMCLKI,
	input USRMCLKTS
);

endmodule
